module hello();

endmodule // hello
